module design;
        initial begin
                $display ("Hello world");
endmodule;
